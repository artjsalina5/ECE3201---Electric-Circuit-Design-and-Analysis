********Problem: P13_66 (b),(c),(d) ***************
******* Main circuit begins here**************
V_CC         VCC 0 10Vdc
Q3         VC12 VC12 VEE Q2N3904
Q1         VC12 IN- VE12 Q2N3906
RL         0 VO  {RL}
I1         VCC VE12 DC 0.1mAdc
Q4         VC24 VC12 VEE Q2N3904
C         VC24 VB7  {Cc}
Q2         VC24 IN+ VE12 Q2N3906
Q6         VO VC24 VEE Q2N3904
Q5         VB7 VC24 VEE Q2N3904
I2         VCC VB7 DC 1mAdc
Q7         VCC VB7 VO Q2N3904
V_EE         0 VEE 10Vdc
V1         IN+ 0  AC 1
+SIN -15.43m 10m 1k 0 0 0
V2         IN- 0  AC -1
+SIN 0 10m 1k 0 0 0
.PARAM  cc=10n rl=5k
******* Main circuit ends here***************

***************** Q2N3906 model begins here ******************************
.model Q2N3906	PNP(Is=1.41f Xti=3 Eg=1.11 Vaf=10000 Bf=100 Ne=1.5 Ise=0
+		Ikf=80m Xtb=1.5 Br=4.977 Nc=2 Isc=0 Ikr=0 Rc=2.5 Cjc=9.728p
+		Mjc=.5776 Vjc=.7 Fc=.5 Cje=8.063p Mje=.3677 Vje=.7 Tr=33.42n
+		Tf=179.3p Itf=.4 Vtf=4 Xtf=6 Rb=10)
***************** Q2N3906 model ends here ******************************

***************** Q2N3904 model begins here ******************************
.model Q2N3904	NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=10000 Bf=100 Ne=1.259
+		Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+		Cjc=3.638p Mjc=.3085 Vjc=.7 Fc=.5 Cje=4.493p Mje=.2593 Vje=.7
+		Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
***************** Q2N3904 model ends here ******************************
******** Analysis begins here****************
.AC  DEC   20  1 1K
*.STEP LIN PARAM cc 0.1n 0.3n 0.025n
.PROBE
.END
******** Analysis ends here****************

