********Example S 16.1 ***************
******* Main circuit begins here**************
V_Vin         IN 0
+PULSE 0 {VDD} 2n 1p 1p 6n 12n
M_M1         OUT IN VDD VDD PMOS0P5
+ L=0.5u
+ W=1.25u
+ AD=1.72E-12
+ AS=1.72E-12
+ PD=5.25e-6
+ PS=5.25E-6
+ M={MP}
C_C10         0 OUT  {CL}
M_M2         OUT IN 0 0 NMOS0P5
+ L=0.5u
+ W=1.25u
+ AD=1.72E-12
+ AS=1.72E-12
+ PD=5.25E-6
+ PS=5.25E-6
+ M={MN}
V_Vsupply         VDD 0 {VDD}
.PARAM  cl=0.5p vdd=3.3 mp=1 mn=1
******* Main circuit ends here**************

************Model for NMOS in 0.5um CMOS Technology begins here*****************
* 		(created by Anas Hamoui & Olivier Trescases)
.model NMOS0P5	NMOS(Level=1 VTO=0.7 GAMMA=0.5 PHI=0.8
+		LD=0.08E-06 WD=0 UO=460 LAMBDA=0.1 TOX=9.5E-9 PB=0.9 CJ=0.57E-3
+		CJSW=120E-12 MJ=0.5 MJSW=0.4 CGDO=0.4E-9 JS=10E-9 CGBO=0.38E-9
+		CGSO=0.4E-9)
************Model for NMOS in 0.5um CMOS Technology ends here*****************

************Model for PMOS in 0.5um CMOS Technology begins here*****************
* 		(created by Anas Hamoui & Olivier Trescases)
.model PMOS0P5	PMOS(Level=1 VTO=-0.8 GAMMA=0.45 PHI=0.8
+		LD=0.09E-06 WD=0 UO=115 LAMBDA=0.2 TOX=9.5E-9 PB=0.9 CJ=0.93E-3
+		CJSW=170E-12 MJ=0.5 MJSW=0.35 CGDO=0.35E-9 JS=5E-9 CGBO=0.38E-9
+		CGSO=0.35E-9)
************Model for PMOS in 0.5um CMOS Technology ends here*****************

******** Analysis begins here****************
.DC [LIN] V_Vin  0 3.3 10m
*.TRAN 	0.01nS  14nS
.PROBE
.END
******** Analysis ends here****************




 
