********Example S 11.2 (Av) ***********************
******* Main circuit begins here**************
V_V4         VIN 0  AC 1Vac
+SIN 0 1m 1k 0 0 0
M_M1         VD1 VIN VD5 0 NMOS4  
+ L=0.2u  
+ W=0.48u  
+ AD=1.72E-12  
+ AS=1.72E-12  
+ PD=5.25E-6  
+ PS=5.25E-6      
+ M=7
M_M3         VD1 VD1 VDD VDD PMOS4  
+ L=0.2u  
+ W=0.64u  
+ AD=1.72E-12  
+ AS=1.72E-12  
+ PD=5.25e-6  
+ PS=5.25E-6      
+ M=15
I_I1         VDD VG5 DC 200uAdc  
M_M5         VD5 VG5 VSS 0 NMOS4  
+ L=0.2u  
+ W=0.48u  
+ AD=1.72E-12  
+ AS=1.72E-12  
+ PD=5.25E-6  
+ PS=5.25E-6      
+ M=14
M_M8         VG5 VG5 VSS 0 NMOS4  
+ L=0.2u  
+ W=0.48u  
+ AD=1.72E-12  
+ AS=1.72E-12  
+ PD=5.25E-6  
+ PS=5.25E-6      
+ M=14
V_V2         0 VSS 1Vdc
M_M4         VD2 VD1 VDD VDD PMOS4  
+ L=0.2u  
+ W=0.64u  
+ AD=1.72E-12  
+ AS=1.72E-12  
+ PD=5.25e-6  
+ PS=5.25E-6      
+ M=15
M_M7         VOUT VG5 VSS 0 NMOS4  
+ L=0.2u  
+ W=0.48u  
+ AD=1.72E-12  
+ AS=1.72E-12  
+ PD=5.25E-6  
+ PS=5.25E-6      
+ M=14
M_M2         VD2 0 VD5 0 NMOS4  
+ L=0.2u  
+ W=0.48u  
+ AD=1.72E-12  
+ AS=1.72E-12  
+ PD=5.25E-6  
+ PS=5.25E-6      
+ M=7
V_V3         VDD 0 1Vdc
M_M6         VDD VD2 VOUT 0 NMOS4  
+ L=0.2u  
+ W=0.48u  
+ AD=1.72E-12  
+ AS=1.72E-12  
+ PD=5.25E-6  
+ PS=5.25E-6      
+ M=14
******* Main circuit ends here**************

*****************PMOS and NMOS models begin here*********************
.model NMOS4	NMOS(LEVEL= 1 VTO=0.5 GAMMA= 0.3  PHI=0.84
+ LAMBDA= 0.08
+ RS=    0.0
+ RD=    0.0
+ CBD=   0.0
+ CBS=   0.0
+ IS=    1.0e-14
+ PB=    0.9
+ CGSO=  0.3665e-9
+ CGDO=   0.3665e-9
+ CGBO=   0.38e-9
+ RSH=   0
+ CJ=    1.6e-3
+ MJ=    0.5
+ CJSW=  2.0405e-10
+ MJSW=  0.200379
+ JS=    8.38e-6
+ TOX= 4.08e-09
+ NSS=   0.0
+ TPG=   1.0
+ LD=    10e-9
+ U0 = 291
+ KF=    0.0
+ AF=    1.0
+ FC=    0.5
+ TNOM=  27
+ )

.model PMOS4	PMOS(LEVEL= 1 VTO=-0.5 KP=86.1e-6  GAMMA= 0.3
+ PHI=   0.8
+ LAMBDA= 0.11
+ RS=    0.0
+ RD=    0.0
+ CBD=   0.0
+ CBS=   0.0
+ IS=    1.0e-14
+ PB=    0.9
+ CGSO=  0.3426e-9
+ CGDO=  0.3426e-9
+ CGBO=  0.35e-9
+ RSH=   0
+ CJ=    1.01574e-03
+ MJ=    0.4490538
+ CJSW=  2.0405e-10
+ MJSW=  0.2931001
+ JS=    4e-7
+ NSS=   0.0
+ TPG=   1.0
+ LD=    10e-9
+ KF=    0.0
+ AF=    1.0
+ FC=    0.5
+ TNOM=  27
+ )
*****************PMOS and NMOS models end here*********************


******** Analysis begins here****************
.OP
.AC  DEC   20  1MEG 5G
.PROBE
.END
******** Analysis ends here****************
