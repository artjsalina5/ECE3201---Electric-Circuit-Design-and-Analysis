********Problem: P8_5		***************
******* Main circuit begins here**************
I1         VDD VG DC 25u
V1         N1 0 0.8Vdc
V2         VDD 0 1.8Vdc
M1         VG VG 0 0 NMOS0P18
+ L=0.54u
+ W=1.74u
+ M=1
M2         VO VG 0 0 NMOS0P18
+ L=0.54u
+ W=6.96u
+ M=1
V3         VO N1  AC 1m
+SIN 0 1m 10k 0 0 0
******* Main circuit ends here**********************************************

***************** NMOS model begins here ******************************
.model NMOS0P18	NMOS(Level=1 VTO=0.5 GAMMA=0.3 PHI=0.84
+		LD=0 WD=0 UO=450 LAMBDA=0.4 TOX=4.08E-9 PB=0.9 CJ=1.6E-3
+		CJSW=2.04E-10 MJ=0.5 MJSW=0.2 CGDO=3.67E-10 JS=8.38E-6 CGBO=3.8E-10
+		CGSO=3.67E-10)
***************** NMOS model ends here *****************************************
******** Analysis begins here****************
.OP
*.AC  DEC   20  1 100K
.PROBE
.END
******** Analysis ends here****************
