********Example PS 2.1(b) (i), (ii), (iii)***************
******* Main circuit begins here**************
R1         N1 0  1k
Vin         N2 0 DC 0Vdc AC 1Vac
R2         N1 OUT  100k
X_A1         N2 N1 OUT OPAMP_MACRO
******* Main circuit ends here **************

******* Opamp macro model begins here **************
.SUBCKT OPAMP_MACRO    IN+ IN- OUT
Ro         OUT N3  75
VOS         N4 IN- 1m
Eb         N3 0 N2 0 1
Rb         N2 N1  16MEG
Cb         0 N2  1n
Ed         N1 0 IN+ N4 1E5
Rid         IN+ N4  2MEG
.ENDS
******* Opamp macro model ends here **************

******** Analysis begins here****************
.OP
.AC  DEC   20  0.1 10MEG
.PROBE
.END
******** Analysis ends here****************
