********Problem: P8_82		***************
******* Main circuit begins here**************
M1         VG12 VG12 0 0 NMOS0P18
+ L=0.54u
+ W=2.7u
+ M=1
M2         N14530 VG12 0 0 NMOS0P18
+ L=0.54u
+ W=27u
+ M=1
M3         VOUT VG34 N14530 0 NMOS0P18
+ L=0.54u
+ W=27u
+ M=1
M4         VG34 VG34 VG12 0 NMOS0P18
+ L=0.54u
+ W=2.7u
+ M=1
I1         VDD VG34 DC 20uAdc
V1         VDD 0 1.8Vdc
V2         VOUT 0  AC 1k
+SIN 0.9 1m 1k 0 0 0
******* Main circuit ends here**********************************************


***************** NMOS model (0.18um) begins here ******************************
.model NMOS0P18	NMOS(Level=1 VTO=0.5 GAMMA=0.3 PHI=0.84
+		LD=0 WD=0 UO=450 LAMBDA=0.55 TOX=4.08E-9 PB=0.9 CJ=1.6E-3
+		CJSW=2.04E-10 MJ=0.5 MJSW=0.2 CGDO=3.67E-10 JS=8.38E-6 CGBO=3.8E-10
+		CGSO=3.67E-10)
***************** NMOS model ends here *****************************************


******** Analysis begins here****************
.OP
*.DC [LIN] V2  0.3 1.0 0.05
*.AC  DEC   20  1 100K
.PROBE
.END
******** Analysis ends here****************
