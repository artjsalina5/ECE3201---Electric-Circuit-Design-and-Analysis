******* Problem: P9_57 **********************
******* Main circuit begins here**************
V_DD         VDD 0 2Vdc
RD2         VOUT2 VDD  107k
RSS         0 VS  20k
RD1         VOUT1 VDD  107k
M1         VOUT1 VG1 VS 0 NMOS0P18
+ L=0.5u
+ W=1.3u
+ M=1
M2         VOUT2 VG2 VS 0 NMOS0P18
+ L=0.5u
+ W=1.3u
+ M=1
VID         VG1 VG2  AC 1m
+SIN 0 1m 1k 0 0 0
VCM         VG2 0 0.95Vdc
******* Main circuit ends here***************

***************** NMOS model begins here ******************************
.model NMOS0P18	NMOS(Level=1 VTO=0.4 GAMMA=0.1 PHI=0.84
+		LD=0 WD=0 UO=450 LAMBDA=0.0 TOX=4.08E-9 PB=0.9 CJ=1.6E-3
+		CJSW=2.04E-10 MJ=0.5 MJSW=0.2 CGDO=3.67E-10 JS=8.38E-6 CGBO=3.8E-10
+		CGSO=3.67E-10)
***************** NMOS model ends here *****************************************

******** Analysis begins here****************
.OP
.DC [LIN] VCM  0 1.5 0.1
*.TRAN 0.01mS  2mS
.PROBE
.END
******** Analysis ends here****************
