********Example S 6.1 ***************
******* Main circuit begins here**************
Q1         N111317 N111357 0 Q2N3904
V1         N111317 0 {VCE}
Ibase         0 N111357 DC {ib}  
.PARAM  ib=10u vce=2v
******* Main circuit ends here**************
**************Model for 2N3904 NPN BJT (from Eval library in Pspice) begins here***********
.model Q2N3904	NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+		Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+		Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+		Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
**************Model for 2N3904 NPN BJT (from Eval library in Pspice) ends here***********
******** Analysis begins here****************
.DC [LIN] Ibase  1u 200u 1u
.PROBE 
.END
******** Analysis ends here****************
