********Example S 7.2 ***************
******* Main circuit begins here**************
C2         N1 VB  {CCI}  
R7         0 VB  {RB}  
V5         IN 0 DC 0Vdc AC 1Vac 
Q2         VC VB VE Q2N3904
V7         VSS 0 {VSS}
R4         VC VDD  {RC}  
R9         0 N2  {RCE}  
R8         VSS VE  {RE}  
C1         VC OUT  {CCO}  
C3         N2 VE  {CB}  
R6         0 OUT  {RL}  
R5         IN N1  {Rsig}  
V6         VDD 0 {VDD}
.PARAM  rc=10k cb=10u re2=1 vss=-5 rb=340k re1=6k cco=10u vdd=5 cci=10u rl=10k
+  rsig=10k rx=1 re=6k rce=130
******* Main circuit ends here**************

**************Model for 2N3904 NPN BJT (from Eval library in Pspice) begins here***********
.model Q2N3904	NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+		Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+		Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+		Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
**************Model for 2N3904 NPN BJT (from Eval library in Pspice) ends here***********

******** Analysis begins here****************
.OP
.AC  DEC   20  1 10MEG
.PROBE 
.END
******** Analysis ends here****************

