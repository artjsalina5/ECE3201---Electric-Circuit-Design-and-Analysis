********Example S 4.1 ***************
******* Main circuit begins here**************
D1         3 6 D1N4148 
D2         5 6 D1N4148 
R3         7 4  {Rload}  
Vsin         1 0  
+SIN 0 169 60 0 0 0
C1         4 6  {C}  
R1         7 6  {R}  
X_Z1         4 7 ZENER_DIODE 
R4         4 0  {Risolation}  
R2         2 1  {Rs}  
X_TX1         0 2 3 4 5 TX 
.PARAM  rs=0.5 risolation=100e6 c=520u rload=200 r=191
******* Main circuit ends here **************


******** Model of ZENER DIODE begins here****************
.SUBCKT ZENER_DIODE 1 2
*connections:       | |
*	       andode |
*		cathode
Dforward 1 2 1mA_diode
Dreverse 2 4 ideal_diode
Vz0 4 3 DC 4.9V
Rz 1 3 10
* diode model statements
.model 1mA_diode D (Is=100pA n=1.679)
.model ideal_diode D (Is=100pA n=0.01)
.ends ZENER_DIODE
******** Model of ZENER DIODE ends here****************

******** Model of 1N4148 Diode (from EVAL library in PSpice) begins here****************
.model D1N4148  D(Is=2.682n N=1.836 Rs=.5664 Ikf=44.17m Xti=3 Eg=1.11 Cjo=4p
+               M=.3333 Vj=.5 Fc=.5 Isr=1.565n Nr=2 Bv=100 Ibv=100u Tt=11.54n)
******** Model of 1N4148 Diode (from EVAL library in PSpice) ends here****************

******** Model of Nonlinear Transformer with Center-Tapped Secondary begins here****************
.subckt TX 1 2 3 4 5 Params: 
Lp 2 1 10mH
Ls1 3 4 52uH
Ls2 4 5 52uH
K1 Lp Ls1 0.999
K2 Lp Ls2 0.999
K3 Ls1 Ls2 0.999
.ends TX
******** Model of Nonlinear Transformer with Center-Tapped Secondary ends here****************

******** Analysis begins here****************
.TRAN 	0.1mS  200mS
.PROBE
.END
******** Analysis ends here****************

