********Problem: P7_101	***************
******* Main circuit begins here**************
V_DD         VDD 0 5Vdc
RD         VDD VD  5k
M1         VD VG 0 0 NMOS0P5
+ L=0.8u
+ W=22u
+ M=1
RG         VG VD  10MEG
******* Main circuit ends here*******************************
***************** NMOS model begins here ********************
.model NMOS0P5	NMOS(Level=1 VTO=0.7 GAMMA=0.5 PHI=0.8
+		LD=0 WD=0 UO=500 LAMBDA=0.001 TOX=9.5E-9 PB=0.9 CJ=0.57E-3
+		CJSW=120E-12 MJ=0.5 MJSW=0.4 CGDO=0.4E-9 JS=10E-9 CGBO=0.38E-9
+		CGSO=0.4E-9)
***************** NMOS model ends here **********************

******** Analysis begins here****************
.op
******** Analysis ends here******************
